/*
*  Name         :dsp_nco.v
*  Description  :
*  Origin       :230507
*  EE           :hel
*/
module dsp_nco #(
    
)(
    
);

endmodule
